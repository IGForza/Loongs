module InstructionMemory(
	input      [32 -1:0] Address, 
	output reg [32 -1:0] Instruction
);
	
	always @(*)
		case (Address[9:2])

			// -------- Paste Binary Instruction Below (Inst-q1-1/Inst-q1-2.txt)

8'd0: Instruction <= 32'h201d0400;
8'd1: Instruction <= 32'h8c080010;
8'd2: Instruction <= 32'hac080000;
8'd3: Instruction <= 32'h20040014;
8'd4: Instruction <= 32'h8c050000;
8'd5: Instruction <= 32'h0c10008f;
8'd6: Instruction <= 32'h8c080004;
8'd7: Instruction <= 32'hac080010;
8'd8: Instruction <= 32'h8c0f0000;
8'd9: Instruction <= 32'h200e0001;
8'd10: Instruction <= 32'h200d0014;
8'd11: Instruction <= 32'h3c18ffff;
8'd12: Instruction <= 32'haf380000;
8'd13: Instruction <= 32'h8db80000;
8'd14: Instruction <= 32'h330c000f;
8'd15: Instruction <= 32'h200b0000;
8'd16: Instruction <= 32'h20100000;
8'd17: Instruction <= 32'h1190001e;
8'd18: Instruction <= 32'h22100001;
8'd19: Instruction <= 32'h1190001e;
8'd20: Instruction <= 32'h22100001;
8'd21: Instruction <= 32'h1190001e;
8'd22: Instruction <= 32'h22100001;
8'd23: Instruction <= 32'h1190001e;
8'd24: Instruction <= 32'h22100001;
8'd25: Instruction <= 32'h1190001e;
8'd26: Instruction <= 32'h22100001;
8'd27: Instruction <= 32'h1190001e;
8'd28: Instruction <= 32'h22100001;
8'd29: Instruction <= 32'h1190001e;
8'd30: Instruction <= 32'h22100001;
8'd31: Instruction <= 32'h1190001e;
8'd32: Instruction <= 32'h22100001;
8'd33: Instruction <= 32'h1190001e;
8'd34: Instruction <= 32'h22100001;
8'd35: Instruction <= 32'h1190001e;
8'd36: Instruction <= 32'h22100001;
8'd37: Instruction <= 32'h1190001e;
8'd38: Instruction <= 32'h22100001;
8'd39: Instruction <= 32'h1190001e;
8'd40: Instruction <= 32'h22100001;
8'd41: Instruction <= 32'h1190001e;
8'd42: Instruction <= 32'h22100001;
8'd43: Instruction <= 32'h1190001e;
8'd44: Instruction <= 32'h22100001;
8'd45: Instruction <= 32'h1190001e;
8'd46: Instruction <= 32'h22100001;
8'd47: Instruction <= 32'h1190001e;
8'd48: Instruction <= 32'h2011003f;
8'd49: Instruction <= 32'h0810004f;
8'd50: Instruction <= 32'h20110006;
8'd51: Instruction <= 32'h0810004f;
8'd52: Instruction <= 32'h2011005b;
8'd53: Instruction <= 32'h0810004f;
8'd54: Instruction <= 32'h2011004f;
8'd55: Instruction <= 32'h0810004f;
8'd56: Instruction <= 32'h20110066;
8'd57: Instruction <= 32'h0810004f;
8'd58: Instruction <= 32'h2011006d;
8'd59: Instruction <= 32'h0810004f;
8'd60: Instruction <= 32'h2011007d;
8'd61: Instruction <= 32'h0810004f;
8'd62: Instruction <= 32'h20110007;
8'd63: Instruction <= 32'h0810004f;
8'd64: Instruction <= 32'h2011007f;
8'd65: Instruction <= 32'h0810004f;
8'd66: Instruction <= 32'h2011006f;
8'd67: Instruction <= 32'h0810004f;
8'd68: Instruction <= 32'h20110077;
8'd69: Instruction <= 32'h0810004f;
8'd70: Instruction <= 32'h201100ff;
8'd71: Instruction <= 32'h0810004f;
8'd72: Instruction <= 32'h20110039;
8'd73: Instruction <= 32'h0810004f;
8'd74: Instruction <= 32'h201100bf;
8'd75: Instruction <= 32'h0810004f;
8'd76: Instruction <= 32'h20110079;
8'd77: Instruction <= 32'h0810004f;
8'd78: Instruction <= 32'h20110071;
8'd79: Instruction <= 32'h200a0000;
8'd80: Instruction <= 32'h116a0006;
8'd81: Instruction <= 32'h214a0001;
8'd82: Instruction <= 32'h116a0008;
8'd83: Instruction <= 32'h214a0001;
8'd84: Instruction <= 32'h116a000a;
8'd85: Instruction <= 32'h214a0001;
8'd86: Instruction <= 32'h116a000e;
8'd87: Instruction <= 32'h22320100;
8'd88: Instruction <= 32'h330c00f0;
8'd89: Instruction <= 32'h000c6102;
8'd90: Instruction <= 32'h08100063;
8'd91: Instruction <= 32'h22330200;
8'd92: Instruction <= 32'h330c0f00;
8'd93: Instruction <= 32'h000c6202;
8'd94: Instruction <= 32'h08100063;
8'd95: Instruction <= 32'h22340400;
8'd96: Instruction <= 32'h330cf000;
8'd97: Instruction <= 32'h000c6302;
8'd98: Instruction <= 32'h08100063;
8'd99: Instruction <= 32'h216b0001;
8'd100: Instruction <= 32'h08100010;
8'd101: Instruction <= 32'h22350800;
8'd102: Instruction <= 32'h20160000;
8'd103: Instruction <= 32'h201c00c8;
8'd104: Instruction <= 32'h201b0000;
8'd105: Instruction <= 32'h20172710;
8'd106: Instruction <= 32'h20090000;
8'd107: Instruction <= 32'h137c001c;
8'd108: Instruction <= 32'h237b0001;
8'd109: Instruction <= 32'h201a0000;
8'd110: Instruction <= 32'haf320000;
8'd111: Instruction <= 32'h20160001;
8'd112: Instruction <= 32'h235a0001;
8'd113: Instruction <= 32'h13570001;
8'd114: Instruction <= 32'h0810006e;
8'd115: Instruction <= 32'h237b0001;
8'd116: Instruction <= 32'h201a0000;
8'd117: Instruction <= 32'haf330000;
8'd118: Instruction <= 32'h20160002;
8'd119: Instruction <= 32'h235a0001;
8'd120: Instruction <= 32'h13570001;
8'd121: Instruction <= 32'h08100075;
8'd122: Instruction <= 32'h237b0001;
8'd123: Instruction <= 32'h201a0000;
8'd124: Instruction <= 32'haf340000;
8'd125: Instruction <= 32'h20160003;
8'd126: Instruction <= 32'h235a0001;
8'd127: Instruction <= 32'h13570001;
8'd128: Instruction <= 32'h0810007c;
8'd129: Instruction <= 32'h237b0001;
8'd130: Instruction <= 32'h201a0000;
8'd131: Instruction <= 32'haf350000;
8'd132: Instruction <= 32'h20160000;
8'd133: Instruction <= 32'h235a0001;
8'd134: Instruction <= 32'h1357ffe3;
8'd135: Instruction <= 32'h08100083;
8'd136: Instruction <= 32'h21ad0004;
8'd137: Instruction <= 32'h21ce0001;
8'd138: Instruction <= 32'h01ee082a;
8'd139: Instruction <= 32'h1020ff81;
8'd140: Instruction <= 32'h3c18fffe;
8'd141: Instruction <= 32'haf380000;
8'd142: Instruction <= 32'h0810008e;
8'd143: Instruction <= 32'hafbf0000;
8'd144: Instruction <= 32'h23bdfffc;
8'd145: Instruction <= 32'h20080001;
8'd146: Instruction <= 32'h00054821;
8'd147: Instruction <= 32'hafa80000;
8'd148: Instruction <= 32'hafa9fffc;
8'd149: Instruction <= 32'h23bdfff8;
8'd150: Instruction <= 32'h00082821;
8'd151: Instruction <= 32'h0c1000a7;
8'd152: Instruction <= 32'h00025021;
8'd153: Instruction <= 32'hac0a000c;
8'd154: Instruction <= 32'h00053021;
8'd155: Instruction <= 32'h8c05000c;
8'd156: Instruction <= 32'h0c1000b8;
8'd157: Instruction <= 32'h23bd0008;
8'd158: Instruction <= 32'h8fa80000;
8'd159: Instruction <= 32'h8fa9fffc;
8'd160: Instruction <= 32'h21080001;
8'd161: Instruction <= 32'h0109502a;
8'd162: Instruction <= 32'h214affff;
8'd163: Instruction <= 32'h1140ffef;
8'd164: Instruction <= 32'h23bd0004;
8'd165: Instruction <= 32'h8fbf0000;
8'd166: Instruction <= 32'h03e00008;
8'd167: Instruction <= 32'h00054080;
8'd168: Instruction <= 32'h01044020;
8'd169: Instruction <= 32'h8d090000;
8'd170: Instruction <= 32'h20a8ffff;
8'd171: Instruction <= 32'h8c0a0004;
8'd172: Instruction <= 32'h214a0001;
8'd173: Instruction <= 32'hac0a0004;
8'd174: Instruction <= 32'h00085880;
8'd175: Instruction <= 32'h01645820;
8'd176: Instruction <= 32'h8d6c0000;
8'd177: Instruction <= 32'h012c082a;
8'd178: Instruction <= 32'h10200003;
8'd179: Instruction <= 32'h2108ffff;
8'd180: Instruction <= 32'h0100082a;
8'd181: Instruction <= 32'h1020fff5;
8'd182: Instruction <= 32'h21020001;
8'd183: Instruction <= 32'h03e00008;
8'd184: Instruction <= 32'h00064080;
8'd185: Instruction <= 32'h01044020;
8'd186: Instruction <= 32'h8d090000;
8'd187: Instruction <= 32'h20c8ffff;
8'd188: Instruction <= 32'h00085080;
8'd189: Instruction <= 32'h01445020;
8'd190: Instruction <= 32'h8d4c0000;
8'd191: Instruction <= 32'had4c0004;
8'd192: Instruction <= 32'h2108ffff;
8'd193: Instruction <= 32'h0105082a;
8'd194: Instruction <= 32'h1020fff9;
8'd195: Instruction <= 32'h00055080;
8'd196: Instruction <= 32'h01445020;
8'd197: Instruction <= 32'had490000;
8'd198: Instruction <= 32'h03e00008;



			// -------- Paste Binary Instruction Above
			
			default: Instruction <= 32'h00000000;
		endcase
		
endmodule
